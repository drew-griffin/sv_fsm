//////////////////////////////////////////////////////////////
// tb_findMax.sv - Testbench to verify that the findMax FSM-D works as specified
//
// Author:	Roy Kravitz (roy.kravitz@pdx.edu) 
// Modified by: Drew Seidel (dseidel@pdx.edu) - closing statement modified for ECE 508 Fall 2022
// Description:
// ------------
// Implements a testbench for the findMax problem on Homework #2.  This testbench
// makes use several of the SystemVerilog verification features including classes
// and constrained randomization and assertions.   These verification constructs are not
// synthesizable.
//
// Original testbench provided by Donald Thomas (Solution is in Problem 7.6)
////////////////////////////////////////////////////////////////
module tb_findMax;

// make use of the SystemVerilog C programming interface
// https://stackoverflow.com/questions/33394999/how-can-i-know-my-current-path-in-system-verilog
import "DPI-C" function string getenv(input string env_name);

// inputs and outputs to the findMax FSM-D
logic start, clk, rst, done;
logic [7:0] inputA, maxValue;

bit [7:0] myMax, savedMax;
int errorCnt = 0;

// instantiate the findMax FSM-D
findMax DUT(.*);

initial begin: monitor_outputs
    $monitor($time,, "state=%s, next_state=%s, start=%b, inputA=%h, done=%b, myMax=%h, maxValue=%h",
        DUT.FSM.STATE, DUT.FSM.NEXT_STATE, start, inputA, done, myMax, maxValue);
end: monitor_outputs

initial begin: clock_reset_gen
    rst = 0;
    rst <= 1;
    #1 rst = 0;
    clk = 0;
    forever #5 clk = ~clk;
end: clock_reset_gen

// number generator (uses constrained randomization)
class pktMax;
    rand bit [7:0] howMany;     // number of unsigned numbers in sequence
    rand bit [7:0] item[];      // dynamic array to hold numbers in sequence
    
    constraint N    {howMany inside {[4:20]};};     // sequences of 4 to 20 unsigned numbers
    constraint arraySize {item.size == howMany;}    // one item for each unsigned number in sequence
endclass

pktMax pkt = new;   // instance of the pktMax class.  Will hold random sequences of unsigned numbers

// stimulus generator and checker
initial begin: stimulus
    // TODO: CHANGE THE GREETING MESSAGE
    $display("ECE (System)Verilog workshop Fall 2022: findMax test - Drew Seidel (dseidel@pdx.edu)");
    $display("Sources: %s\n", getenv("PWD"));
    
    start = 0;
    repeat(20) begin: gen_test_cases    // generate/check 20 sequences
        byte i;
        
        @(posedge clk);
        // fill item[] with random numbers for the sequence
        assert(pkt.randomize()) else $error("Problems generating random numbers");
        
        // deliver all the unsigned numbers in the sequence to the DUT and keep track
        // of the maximum number (myMax) which will be compared to the max number generated by the DUT
        // howMany contains is the length of the sequence
        for (i = 0, myMax = 0; i < pkt.howMany; i++) begin: apply_test_case
            inputA <= pkt.item[i];
            myMax <= (pkt.item[i] < myMax) ? myMax : pkt.item[i];
            start <= 1;
            @(posedge clk);
        end: apply_test_case
        start <= 0;
        @(posedge clk);
        savedMax = myMax;
        if (myMax == maxValue) begin
            $display("Correct max (%h) found", maxValue);
        end
        else begin
            $display("Incorrect max (%h) found, should be %h", maxValue, myMax);
            errorCnt++;
        end
            
        if ((pkt.howMany % 8'h03) == 8'h03)
            @(posedge clk);  // start comes back immediately now and then
    end: gen_test_cases
    
    @(posedge clk);
    if (errorCnt == 0)
        $display("Congratulations!  Your implementation passes the testbench");
    else
        $display("Nice try, but you had %d errors...take a break, do some debug, and try again", errorCnt);
        
    $display("End simulation of findMax test - Drew Seidel (dseidel@pdx.edu)\n");
    $stop;
end:  stimulus

endmodule: tb_findMax
    
        
